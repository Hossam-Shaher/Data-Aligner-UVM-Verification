`ifndef ALGN_IF_SV
  `define ALGN_IF_SV

  interface algn_if(input clk);
    	
    logic reset_n;
    
    logic irq;

  endinterface

`endif