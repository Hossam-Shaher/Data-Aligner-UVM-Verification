`ifndef APB_SEQUENCER_SV
  `define APB_SEQUENCER_SV

  typedef class apb_seq_item_drv;

  typedef uvm_sequencer#(apb_seq_item_drv) apb_sequencer; 

`endif //APB_SEQUENCER_SV